module Experiment6(); // 4-bit ALU

//Declaring general variables

logic in [0:14];
logic out [0:12];

int outf,i;

initial begin

//Reading input and state text files

  $readmemb("C:\\Digikitv3.1Win64\\input.txt",in);

//Assigning default values of the output variables

  for(i=0;i<13;i=i+1)
  begin
    out[i] = 1'bz;
  end
end

//TOP MODULE FUNCTIONS

logic [4:0] dutout;
//5-bit final ALU output including the final Carry Flag

logic [3:0] A,B,not4b,and4b,or4b,xor4b,inc4b,dec4b,add4b,sub4b;
// 4-bit Inputs A B and Outputs for 8 ALU Functions

logic Cin,Cout_inc,Cout_dec,Cout_add,Cout_sub,Carry,sel2,sel1,sel0,enbar;
//Carry bits and Function Select bits

Logic_4bit logic_4b(A,B,not4b,and4b,or4b,xor4b);
// 4-bit Inputs and Outputs for Logic Functions

Arithmetic_4bit arith_4b(A,B,Cin,inc4b,dec4b,add4b,sub4b,Cout_inc,Cout_dec,Cout_add,Cout_sub);
// 4-bit Inputs and 5-bit Outputs including Carry for Arithmetic Functions

MUX_4input_1bit MUX4(Cout_inc,Cout_dec,Cout_add,Cout_sub,sel1,sel0,enbar,Carry);
//Carry generated by Arithmetic functions

and C_Flag(dutout[4],sel2,Carry);
// Final Carry flag generated by the ALU

MUX_8input_4bit Mux8(not4b,and4b,or4b,xor4b,inc4b,dec4b,add4b,sub4b,sel2,sel1,sel0,enbar,dutout[3:0]);
//Final 4-bit ALU output selected by the Function select

initial begin

// Assignments of Switches
  A[3] = in[0];
  A[2] = in[1];
  A[1] = in[2];
  A[0] = in[3];
  B[3] = in[4];
  B[2] = in[5];
  B[1] = in[6];
  B[0] = in[7];
   Cin = in[8];
  sel2 = in[11];
  sel1 = in[12];
  sel0 = in[13];
  enbar= in[14];

#5
// Assignments of output variables to LEDs

    for(i=0;i<5;i++)
    begin
      out[i] = dutout[4-i];
    end
end

initial begin
//Generating output text file

  #5 outf = $fopen("C:\\Digikitv3.1Win64\\output.txt","w");
  #5 $fwrite(outf,"output1 %0b output2 %0b output3 %0b output4 %0b output5 %0b output6 %0b output7 %0b output8 %0b output9 %0b output10 %0b output11 %0b output12 %0b output13 %0b",out[0],out[1],out[2],out[3],out[4],out[5],out[6],out[7],out[8],out[9],out[10],out[11],out[12]);
  #5 $fclose(outf);

end
endmodule  //End of Top Module



module Logic_4bit(A,B,not4b,and4b,or4b,xor4b);
  input [3:0] A,B;
  output [4:0] not4b,and4b,or4b,xor4b;

  assign not4b = ~A;
  assign and4b = A & B;
  assign or4b = A | B;
  assign xor4b = A ^ B;
endmodule

module Arithmetic_4bit(A,B,Cin,inc4b,dec4b,add4b,sub4b,Cout_inc,Cout_dec,Cout_add,Cout_sub);
  input [3:0] A,B;
  input Cin;
  output [3:0] inc4b,dec4b,add4b,sub4b;
  output Cout_inc,Cout_dec,Cout_add,Cout_sub;

  assign {Cout_inc, inc4b} = A + 1'b1;
  assign {Cout_dec, dec4b} = A - 1'b1;
  assign {Cout_add, add4b} = A + B + Cin;
  assign {Cout_sub, sub4b} = A - B - Cin;
endmodule

module MUX_4input_1bit(Cout_inc,Cout_dec,Cout_add,Cout_sub,sel1,sel0,enbar,Carry);
  input Cout_inc,Cout_dec,Cout_add,Cout_sub,sel1,sel0,enbar;
  output Carry;

  assign Carry = enbar?1'b0:(sel1?(sel0?Cout_sub:Cout_add):(sel0?Cout_dec:Cout_inc));
endmodule

module MUX_8input_4bit(not4b,and4b,or4b,xor4b,inc4b,dec4b,add4b,sub4b,sel2,sel1,sel0,enbar,dutout[3:0]);
  input [3:0] not4b,and4b,or4b,xor4b,inc4b,dec4b,add4b,sub4b;
  input sel2,sel1,sel0,enbar;
  output [3:0] dutout;

  assign dutout = enbar?4'b0:(sel2?(sel1?(sel0?sub4b:add4b):(sel0?dec4b:inc4b)):(sel1?(sel0?xor4b:or4b):(sel0?and4b:not4b)));
endmodule
